///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: CPU_MultiCycle (CLK=100)
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// Extended By: CDA3102 students
// License: MIT, (C) 2020-2023 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbenchLui();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Inputs: clk, reset (1-bit)
   reg clk, rst;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Outputs: PC (32-bit), OPCODE (6-bit), FUNCTCODE (6-bit), STATE (5-bit)
wire[31:0] PC;
wire[31:26] OPCODE;
wire[31:26] FUNCTCODE;
wire[4:0] STATE;
///////////////////////////////////////////////////////////////////////////////////

   integer address;

///////////////////////////////////////////////////////////////////////////////////
// Component is CLOCKED
// Set clk period to 100 in wave
// Approximating clock period as 100 (one access to RAM)
localparam CLK_PERIOD=100;
///////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////////////
// CPU will perform check once PC hits this value
// Note for this CPU you want to go *two* past the end
// Because PC=PC+4 when the instruction is still running, in state 0
localparam TERMINALPC=12;
////////////////////////////////////////////////////////////////////////////////////////////////////

   CPU_MultiCycle myCPU(.clk(clk), .reset(rst), ._PC(PC), .FUNCTCODE(FUNCTCODE), .OPCODE(OPCODE), .state(STATE));
   
   initial begin
     ////////////////////////////////////////////////////////////////////////////////////////////////////////////
      // Initialize Instruction Memory with MIPS Bubble Sort         //          INSTRUCTION                    PC
      myCPU.b2v_IDM.memory[0] = 'b00111100000010000000000000000001;  //          lui $t0, 1 	 		0	
      myCPU.b2v_IDM.memory[1] = 'b00110101000010000000000000000011;  //          ori $t0, $t0, 3 		1	
      ////////////////////////////////////////////////////////////////////////////////////////////////////////////

      /////////////////////////////////////////////////////////////////////////////////////////////
      // Turn power on for 1 tick
      rst <= 1;  # (CLK_PERIOD);
      /////////////////////////////////////////////////////////////////////////////////////////////
      rst <= 0; 
   end


  always@(posedge clk)
    begin
        ///////////////////////////////////////////////////////////////////////////////////
        if(PC === TERMINALPC) begin
          $display("Testing lui with immediate=1 and ori with immediate=3");
          verifyEqual32(myCPU.b2v_myRF.contents_t0, 65539);
          $display("CPU functional");
          $stop;
         end
        ///////////////////////////////////////////////////////////////////////////////////
   end
 
endmodule
