///////////////////////////////////////////////////////////////////////////////////
// Component: MicroROM
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// Extended By: CDA3102 students
// License: MIT, (C) 2020-2022 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module MicroROM(state, microinstruction);
///////////////////////////////////////////////////////////////////////////////////
// Input: state (4-bit)
  input [4:0] state; 
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Output: microinstruction (18-bit)
  output wire [17:0] microinstruction;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Internal: ROM
  reg [17:0] ROM[15:0];
///////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////
  // PUT MICROINSTRUCTIONS HERE
  // Bit Order: PCWrite, PCWriteCond, IorD, MemWrite, IRWrite, MemToReg (2),
  //            PCSrc (2), ALUOp (2), ALUSrcB (2), ALUSrcA, RegWrite,
  //            RegDst, isBNE, LOWrite
  //////////////////////////////////////////////////////////////////////
  initial begin
  ROM[5'b00000] = 		18'b100010000000100000;	// State 0
  ROM[5'b00001] =		18'b000000000001100000;	// State 1
  ROM[5'b00010] =		18'b000000000001010000;	// State 2
  ROM[5'b00011] =		18'b001000000000000000; // State 3
  ROM[5'b00100] =		18'b000000100000001000;	// State 4
  ROM[5'b00101] =		18'b001100000000000000;	// State 5
  ROM[5'b00110] =		18'b000000000100010000; // State 6
  ROM[5'b00111] = 		18'b000000000000001100; // State 7
  ROM[5'b01000] = 		18'b010000001010010000;	// State 8
  ROM[5'b01001] = 		18'b100000010000000000;	// State 9
  ROM[5'b01010] =	     	18'b000000000000001000;	// State 10
  ROM[5'b01011] =                18'b010000001010010010; // State 11
  ROM[5'b01100] =                18'b000000000111010000; // State 12  
  ROM[5'b01101] =                18'b000000000000000001; // State 13
  ROM[5'b01110] =                18'b000001000000001100; // State 14
  ////////////////////////////////////////////////////////////////////////
  end

  ////////////////////////////////////////////////////////////////////////
  // Microinstruction stored in ROM, address is the state
  assign microinstruction = ROM[state];
  ////////////////////////////////////////////////////////////////////////

endmodule
