///////////////////////////////////////////////////////////////////////////////////
// Component: MicroROM
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// Extended By: CDA3102 students
// License: MIT, (C) 2020-2022 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module MicroROM(state, microinstruction);
///////////////////////////////////////////////////////////////////////////////////
// Input: state (4-bit)
  input [3:0] state; 
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Output: microinstruction (17-bit)
  output wire [16:0] microinstruction;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Internal: ROM
  reg [16:0] ROM[15:0];
///////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////
  // PUT MICROINSTRUCTIONS HERE
  // Bit Order: PCWrite, PCWriteCond, IorD, MemWrite, IRWrite, MemToReg,
  //            PCSrc (2), ALUOp (2), ALUSrcB (2), ALUSrcA, RegWrite,
  //            RegDst, isBNE, AddrCtl
  //////////////////////////////////////////////////////////////////////
  initial begin
  ROM[4'b0000] = 		17'b10001000000100001;	// State 0
  ROM[4'b0001] =		17'b00000000001100000;	// State 1
  ROM[4'b0010] =		17'b00000000001010000;	// State 2
  ROM[4'b0011] =		17'b00100000000000001; 	// State 3
  ROM[4'b0100] =		17'b00000100000001000;	// State 4
  ROM[4'b0101] =		17'b00110000000000000;	// State 5
  ROM[4'b0110] =		17'b00000000100010001; 	// State 6
  ROM[4'b0111] = 		17'b00000000000001100; 	// State 7
  ROM[4'b1000] = 		17'b01000001010010000;	// State 8
  ROM[4'b1001] = 		17'b10000010000000000;	// State 9
  ROM[4'b1010] =  		17'b00000000001010001;	// State 10
  ROM[4'b1011] =	     	17'b00000000000001000;	// State 11
  ROM[4'b1100] =                17'b01000001010010010;  // State 12
  ROM[4'b1101] =                17'b00000000111010000;  // State 13  
  ////////////////////////////////////////////////////////////////////////
  end

  ////////////////////////////////////////////////////////////////////////
  // Microinstruction stored in ROM, address is the state
  assign microinstruction = ROM[state];
  ////////////////////////////////////////////////////////////////////////

endmodule
